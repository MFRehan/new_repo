module top()


endmodule
